CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
50 0 30 90 10
175 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
343 176 456 273
9437202 0
0
6 Title:
5 Name:
0
0
0
68
14 Logic Display~
6 1389 152 0 1 2
10 23
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3679 0 0
2
44470.6 3
0
14 Logic Display~
6 1406 152 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9342 0 0
2
44470.6 2
0
14 Logic Display~
6 1439 151 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3623 0 0
2
44470.6 1
0
14 Logic Display~
6 1422 151 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3722 0 0
2
44470.6 0
0
13 Quad 3-State~
48 1399 219 0 9 19
0 26 25 24 23 73 74 75 76 32
0
0 0 4704 602
8 QUAD3STA
-28 -44 28 -36
3 U18
42 -2 63 6
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 512 1 0 0 0
1 U
8993 0 0
2
44470.6 0
0
13 Logic Switch~
5 820 123 0 1 11
0 5
0
0 0 20592 0
2 0V
-6 -16 8 -8
3 V33
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3723 0 0
2
44470.6 0
0
13 Logic Switch~
5 822 168 0 1 11
0 3
0
0 0 20592 0
2 0V
-6 -16 8 -8
3 V32
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6244 0 0
2
44470.6 3
0
13 Logic Switch~
5 822 144 0 1 11
0 4
0
0 0 20592 0
2 0V
-6 -16 8 -8
3 V31
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6421 0 0
2
44470.6 2
0
13 Logic Switch~
5 823 191 0 1 11
0 2
0
0 0 20592 0
2 0V
-6 -16 8 -8
3 V30
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7743 0 0
2
44470.6 1
0
13 Logic Switch~
5 823 212 0 1 11
0 6
0
0 0 20592 0
2 0V
-6 -16 8 -8
3 V29
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9840 0 0
2
44470.6 0
0
13 Logic Switch~
5 1099 444 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 20592 270
2 5V
-6 -16 8 -8
3 V28
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6910 0 0
2
44470.6 0
0
13 Logic Switch~
5 522 444 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 20592 270
2 5V
-6 -16 8 -8
3 V27
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
449 0 0
2
44470.6 0
0
13 Logic Switch~
5 131 438 0 1 11
0 9
0
0 0 20592 0
2 0V
-6 -16 8 -8
3 V26
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8761 0 0
2
44470.6 0
0
13 Logic Switch~
5 132 484 0 1 11
0 52
0
0 0 20592 0
2 0V
-6 -16 8 -8
3 V25
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6748 0 0
2
44470.5 38
0
13 Logic Switch~
5 131 468 0 1 11
0 37
0
0 0 20592 0
2 0V
-6 -16 8 -8
3 V24
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7393 0 0
2
44470.5 37
0
13 Logic Switch~
5 130 452 0 1 11
0 34
0
0 0 20592 0
2 0V
-6 -16 8 -8
3 V23
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7699 0 0
2
44470.5 36
0
13 Logic Switch~
5 142 172 0 1 11
0 30
0
0 0 20592 0
2 0V
-6 -16 8 -8
3 V22
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6638 0 0
2
44470.5 35
0
13 Logic Switch~
5 141 152 0 1 11
0 29
0
0 0 20592 0
2 0V
-6 -16 8 -8
3 V21
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4595 0 0
2
44470.5 34
0
13 Logic Switch~
5 141 114 0 1 11
0 31
0
0 0 20592 0
2 0V
-6 -16 8 -8
3 V20
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9395 0 0
2
44470.5 33
0
13 Logic Switch~
5 143 133 0 10 11
0 28 0 0 0 0 0 0 0 0
1
0
0 0 20592 0
2 5V
-6 -16 8 -8
3 V17
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3303 0 0
2
44470.5 32
0
13 Logic Switch~
5 134 382 0 1 11
0 27
0
0 0 20592 0
2 0V
-6 -16 8 -8
3 V19
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4498 0 0
2
44470.5 31
0
13 Logic Switch~
5 133 400 0 1 11
0 57
0
0 0 20592 0
2 0V
-6 -16 8 -8
3 V18
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9728 0 0
2
44470.5 30
0
13 Logic Switch~
5 134 416 0 10 11
0 39 0 0 0 0 0 0 0 0
1
0
0 0 20592 0
2 5V
-6 -16 8 -8
3 V16
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3789 0 0
2
44470.5 29
0
13 Logic Switch~
5 135 349 0 1 11
0 41
0
0 0 20592 0
2 0V
-6 -16 8 -8
3 V15
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3978 0 0
2
44470.5 28
0
13 Logic Switch~
5 134 366 0 1 11
0 40
0
0 0 20592 0
2 0V
-6 -16 8 -8
3 V14
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3494 0 0
2
44470.5 27
0
13 Logic Switch~
5 134 333 0 1 11
0 42
0
0 0 20592 0
2 0V
-6 -16 8 -8
3 V13
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3507 0 0
2
44470.5 26
0
13 Logic Switch~
5 135 315 0 1 11
0 43
0
0 0 20592 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5151 0 0
2
44470.5 25
0
5 4069~
219 1223 242 0 2 22
0 9 10
0
0 0 624 90
4 4069
-7 -24 21 -16
4 U17E
17 -2 45 6
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 5 4 0
1 U
3701 0 0
2
44470.6 0
0
14 Logic Display~
6 1215 470 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L20
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8585 0 0
2
44470.6 3
0
14 Logic Display~
6 1232 470 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8809 0 0
2
44470.6 2
0
14 Logic Display~
6 1199 471 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5993 0 0
2
44470.6 1
0
14 Logic Display~
6 1182 471 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8654 0 0
2
44470.6 0
0
14 Logic Display~
6 633 469 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7223 0 0
2
44470.6 3
0
14 Logic Display~
6 650 469 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3641 0 0
2
44470.6 2
0
14 Logic Display~
6 617 470 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3104 0 0
2
44470.6 1
0
14 Logic Display~
6 600 470 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3296 0 0
2
44470.6 0
0
14 Logic Display~
6 989 99 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8534 0 0
2
44470.5 3
0
14 Logic Display~
6 1006 99 0 1 2
10 20
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
949 0 0
2
44470.5 2
0
14 Logic Display~
6 1039 98 0 1 2
10 22
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3371 0 0
2
44470.5 1
0
14 Logic Display~
6 1022 98 0 1 2
10 21
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7311 0 0
2
44470.5 0
0
14 Logic Display~
6 541 196 0 1 2
10 25
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3409 0 0
2
44470.5 1
0
14 Logic Display~
6 558 196 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3526 0 0
2
44470.5 0
0
14 Logic Display~
6 525 197 0 1 2
10 24
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4129 0 0
2
44470.5 0
0
14 Logic Display~
6 508 197 0 1 2
10 23
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6278 0 0
2
44470.5 0
0
5 4069~
219 1318 242 0 2 22
0 57 32
0
0 0 624 90
4 4069
-7 -24 21 -16
4 U17D
17 -2 45 6
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 4 4 0
1 U
3482 0 0
2
44470.5 24
0
5 4069~
219 278 274 0 2 22
0 27 33
0
0 0 624 90
4 4069
-7 -24 21 -16
4 U17C
17 -2 45 6
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 3 4 0
1 U
8323 0 0
2
44470.5 23
0
5 4069~
219 1045 243 0 2 22
0 34 35
0
0 0 624 90
4 4069
-7 -24 21 -16
4 U17B
17 -2 45 6
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 2 4 0
1 U
3984 0 0
2
44470.5 21
0
13 Quad 3-State~
48 1087 222 0 9 19
0 19 20 21 22 23 24 25 26 35
0
0 0 4720 270
8 QUAD3STA
-28 -44 28 -36
3 U16
1 -1 22 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
7622 0 0
2
44470.5 20
0
5 4069~
219 956 237 0 2 22
0 37 36
0
0 0 624 90
4 4069
-7 -24 21 -16
4 U17A
17 -2 45 6
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 1 4 0
1 U
816 0 0
2
44470.5 19
0
13 Quad 3-State~
48 1183 221 0 9 19
0 26 25 24 23 22 21 20 19 10
0
0 0 4720 90
8 QUAD3STA
-28 -44 28 -36
2 U2
-23 -1 -9 7
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
4656 0 0
2
44470.5 18
0
5 4069~
219 1293 449 0 2 22
0 40 47
0
0 0 624 270
4 4069
-7 -24 21 -16
4 U15F
17 -8 45 0
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 6 3 0
1 U
6356 0 0
2
44470.5 17
0
5 4069~
219 848 464 0 2 22
0 39 46
0
0 0 624 270
4 4069
-7 -24 21 -16
4 U15E
17 -8 45 0
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
7479 0 0
2
44470.5 16
0
5 4069~
219 715 452 0 2 22
0 41 38
0
0 0 624 270
4 4069
-7 -24 21 -16
4 U15D
17 -8 45 0
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
5690 0 0
2
44470.5 15
0
13 Quad 3-State~
48 1296 525 0 9 19
0 26 25 24 23 14 13 12 11 47
0
0 0 4720 180
8 QUAD3STA
-28 -44 28 -36
3 U10
-10 46 11 54
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
5617 0 0
2
44470.5 14
0
13 Quad 3-State~
48 718 526 0 9 19
0 18 17 16 15 26 25 24 23 38
0
0 0 4720 692
8 QUAD3STA
-28 -44 28 -36
2 U4
-7 46 7 54
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
3903 0 0
2
44470.5 13
0
13 Quad 3-State~
48 889 501 0 9 19
0 51 49 48 50 26 25 24 23 46
0
0 0 4720 602
8 QUAD3STA
-28 -44 28 -36
3 U14
42 -2 63 6
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
4452 0 0
2
44470.5 12
0
5 4030~
219 1049 737 0 3 22
0 52 12 54
0
0 0 624 180
4 4030
-7 -24 21 -16
4 U13D
-5 -25 23 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
6282 0 0
2
44470.5 11
0
5 4030~
219 1050 770 0 3 22
0 52 11 53
0
0 0 624 180
4 4030
-7 -24 21 -16
4 U13C
-5 -25 23 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
7187 0 0
2
44470.5 10
0
5 4030~
219 1050 701 0 3 22
0 52 13 55
0
0 0 624 180
4 4030
-7 -24 21 -16
4 U13B
-5 -25 23 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
6866 0 0
2
44470.5 9
0
5 4030~
219 1049 668 0 3 22
0 52 14 56
0
0 0 624 180
4 4030
-7 -24 21 -16
4 U13A
-5 -25 23 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
7670 0 0
2
44470.5 8
0
7 74LS283
152 901 615 0 14 29
0 15 16 17 18 53 54 55 56 52
50 48 49 51 77
0
0 0 4848 90
6 74F283
-21 -60 21 -52
3 U12
56 -3 77 5
0
15 DVCC=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 14 3 5 11 15 2 6 7
10 13 1 4 9 12 14 3 5 11
15 2 6 7 10 13 1 4 9 0
65 0 0 512 0 0 0 0
1 U
951 0 0
2
44470.5 7
0
7 74LS273
150 1136 512 0 18 37
0 7 44 78 79 80 81 23 24 25
26 82 83 84 85 11 12 13 14
0
0 0 4848 0
6 74F273
-21 -60 21 -52
3 U11
-10 -61 11 -53
0
16 DVCC=20;DGND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 0 0 0 0
1 U
9536 0 0
2
44470.5 6
0
5 4081~
219 1068 443 0 3 22
0 37 42 44
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U9B
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
5495 0 0
2
44470.5 5
0
5 4081~
219 491 453 0 3 22
0 37 43 45
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U9A
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
8152 0 0
2
44470.5 4
0
4 4505
219 144 630 0 12 25
0 86 87 88 89 90 91 92 93 94
95 96 97
0
0 0 4848 0
4 4505
-14 -60 14 -52
2 U8
-7 -61 7 -53
0
15 DVDD=14;DGND=7;
126 %D [%14bi %7bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %12i]
+ [%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %12o %11o] %M
0
12 type:digital
5 DIP14
25

0 12 11 4 3 2 1 5 6 8
9 10 13 12 11 4 3 2 1 5
6 8 9 10 13 0
65 0 0 512 0 0 0 0
1 U
6223 0 0
2
44470.5 3
0
6 1K RAM
79 906 141 0 20 41
0 98 99 100 101 102 5 4 3 2
6 103 104 105 106 19 20 21 22 36
34
0
0 0 4848 0
5 RAM1K
-17 -19 18 -11
2 U7
-7 -70 7 -62
0
16 DVCC=22;DGND=11;
214 %D [%22bi %11bi  %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i %13i %14i %15i %16i %17i %18i %19i %20i]
+ [%22bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o  %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o] %M
0
12 type:digital
5 DIP22
41

0 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 1 2 3 4 5 6 7 8 9
10 12 13 14 15 16 17 18 19 20
21 0
65 0 0 512 0 0 0 0
1 U
5441 0 0
2
44470.5 2
0
7 74LS273
150 559 513 0 18 37
0 8 45 107 108 109 110 23 24 25
26 111 112 113 114 15 16 17 18
0
0 0 4848 0
6 74F273
-21 -60 21 -52
2 U3
-7 -61 7 -53
0
16 DVCC=20;DGND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 512 0 0 0 0
1 U
3189 0 0
2
44470.5 1
0
13 Quad 3-State~
48 254 210 0 9 19
0 30 29 28 31 26 25 24 23 33
0
0 0 4720 0
8 QUAD3STA
-28 -44 28 -36
2 U1
-7 -46 7 -38
0
15 DVCC=16;DGND=8;
85 %D [%16bi %8bi %1i %2i %3i %4i %9i]
+ [%16bo %1o %2o %3o %4o %9o %5o %6o %7o %8o] %M
0
12 type:digital
5 DIP16
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
65 0 0 0 1 0 0 0
1 U
8460 0 0
2
44470.5 0
0
138
1 5 0 0 0 0 0 3 5 0 0 3
1439 169
1439 198
1432 198
6 1 0 0 0 16 0 5 4 0 0 3
1420 198
1420 169
1422 169
1 7 0 0 0 0 0 2 5 0 0 3
1406 170
1408 170
1408 198
1 8 0 0 0 0 0 1 5 0 0 3
1389 170
1389 198
1396 198
2 9 0 0 0 0 0 45 5 0 0 3
1321 224
1321 222
1360 222
1 0 0 0 0 0 0 45 0 0 121 2
1321 260
1321 342
0 1 0 0 0 8320 0 0 22 0 0 4
1480 336
246 336
246 400
145 400
9 1 2 0 0 12416 0 66 9 0 0 4
874 177
857 177
857 191
835 191
1 8 3 0 0 4224 0 7 66 0 0 2
834 168
874 168
1 7 4 0 0 8320 0 8 66 0 0 5
834 144
834 145
857 145
857 159
874 159
1 6 5 0 0 4224 0 6 66 0 0 4
832 123
864 123
864 150
874 150
1 10 6 0 0 4224 0 10 66 0 0 4
835 212
863 212
863 186
874 186
1 1 7 0 0 4224 0 11 62 0 0 3
1099 456
1099 476
1098 476
1 1 8 0 0 8320 0 12 67 0 0 3
522 456
521 456
521 477
1 0 9 0 0 4096 0 28 0 0 18 2
1226 260
1226 353
9 2 10 0 0 4224 0 50 28 0 0 2
1222 224
1226 224
1 0 9 0 0 0 0 13 0 0 18 3
143 438
143 440
139 440
1 0 9 0 0 12416 0 0 0 0 0 4
131 440
270 440
270 353
1467 353
1 0 11 0 0 4096 0 32 0 0 107 2
1182 489
1182 530
1 0 12 0 0 4096 0 31 0 0 108 2
1199 489
1199 539
1 0 13 0 0 4096 0 29 0 0 109 2
1215 488
1215 548
1 0 14 0 0 4096 0 30 0 0 110 2
1232 488
1232 557
1 0 15 0 0 4096 0 36 0 0 127 2
600 488
600 531
1 0 16 0 0 4096 0 35 0 0 128 2
617 488
617 540
1 0 17 0 0 4096 0 33 0 0 129 2
633 487
633 549
1 0 18 0 0 4096 0 34 0 0 130 2
650 487
650 558
1 0 19 0 0 4096 0 37 0 0 63 2
989 117
989 159
1 0 20 0 0 4096 0 38 0 0 64 2
1006 117
1006 168
1 0 21 0 0 4096 0 40 0 0 65 2
1022 116
1022 177
1 0 22 0 0 4096 0 39 0 0 66 2
1039 116
1039 186
1 0 23 0 0 4096 0 44 0 0 135 2
508 215
508 283
1 0 24 0 0 4096 0 43 0 0 136 2
525 215
525 277
1 0 25 0 0 4096 0 41 0 0 137 2
541 214
541 271
1 0 26 0 0 4096 0 42 0 0 138 2
558 214
558 265
1 0 27 0 0 4096 0 46 0 0 122 2
281 292
281 330
1 3 28 0 0 12416 0 20 68 0 0 5
155 133
155 132
178 132
178 204
230 204
1 2 29 0 0 12416 0 18 68 0 0 4
153 152
167 152
167 192
230 192
1 1 30 0 0 8320 0 17 68 0 0 3
154 172
154 180
230 180
1 4 31 0 0 8320 0 19 68 0 0 4
153 114
190 114
190 216
230 216
2 9 33 0 0 8320 0 46 68 0 0 4
281 256
281 250
254 250
254 252
20 0 34 0 0 8192 0 66 0 0 52 3
944 114
945 114
945 361
1 0 34 0 0 0 0 47 0 0 52 2
1048 261
1048 361
2 9 35 0 0 0 0 47 48 0 0 2
1048 225
1048 225
1 0 19 0 0 0 0 48 0 0 63 2
1120 201
1120 159
2 0 20 0 0 0 0 48 0 0 64 2
1108 201
1108 168
3 0 21 0 0 0 0 48 0 0 65 2
1096 201
1096 177
4 0 22 0 0 0 0 48 0 0 66 2
1084 201
1084 186
5 0 23 0 0 0 0 48 0 0 135 2
1120 249
1120 283
6 0 24 0 0 0 0 48 0 0 136 2
1108 249
1108 277
7 0 25 0 0 0 0 48 0 0 137 2
1096 249
1096 271
8 0 26 0 0 0 0 48 0 0 138 2
1084 249
1084 265
1 0 34 0 0 12416 0 16 0 0 0 4
142 452
281 452
281 361
1478 361
2 19 36 0 0 4224 0 49 66 0 0 3
959 219
959 105
944 105
1 0 37 0 0 4096 0 49 0 0 116 2
959 255
959 369
8 0 19 0 0 0 0 50 0 0 63 2
1186 200
1186 159
7 0 20 0 0 0 0 50 0 0 64 2
1174 200
1174 168
6 0 21 0 0 0 0 50 0 0 65 2
1162 200
1162 177
5 0 22 0 0 0 0 50 0 0 66 2
1150 200
1150 186
4 0 23 0 0 0 0 50 0 0 135 2
1186 248
1186 283
3 0 24 0 0 0 0 50 0 0 136 2
1174 248
1174 277
2 0 25 0 0 0 0 50 0 0 137 2
1162 248
1162 271
1 0 26 0 0 0 0 50 0 0 138 2
1150 248
1150 265
15 0 19 0 0 4224 0 66 0 0 0 2
938 159
1279 159
16 0 20 0 0 4224 0 66 0 0 0 2
938 168
1278 168
17 0 21 0 0 4224 0 66 0 0 0 2
938 177
1279 177
18 0 22 0 0 4224 0 66 0 0 0 2
938 186
1278 186
2 9 38 0 0 4224 0 53 55 0 0 2
718 470
718 490
1 0 39 0 0 4096 0 52 0 0 121 2
851 446
851 342
1 0 40 0 0 4096 0 51 0 0 123 2
1296 431
1296 324
1 0 41 0 0 4096 0 53 0 0 124 2
718 434
718 318
2 0 42 0 0 4096 0 63 0 0 125 2
1057 421
1057 311
2 0 43 0 0 4096 0 64 0 0 126 2
480 431
480 305
3 2 44 0 0 8320 0 63 62 0 0 3
1066 466
1066 485
1104 485
2 3 45 0 0 4224 0 67 64 0 0 3
527 486
489 486
489 476
2 9 46 0 0 4224 0 52 56 0 0 3
851 482
851 504
850 504
2 9 47 0 0 4224 0 51 54 0 0 2
1296 467
1296 489
8 0 23 0 0 4096 0 56 0 0 135 2
886 480
886 283
7 0 24 0 0 4096 0 56 0 0 136 2
898 480
898 277
6 0 25 0 0 4096 0 56 0 0 137 2
910 480
910 271
5 0 26 0 0 4096 0 56 0 0 138 2
922 480
922 265
11 3 48 0 0 8320 0 61 56 0 0 3
899 585
898 585
898 528
12 2 49 0 0 12416 0 61 56 0 0 4
908 585
908 576
910 576
910 528
10 4 50 0 0 12416 0 61 56 0 0 4
890 585
890 580
886 580
886 528
13 1 51 0 0 12416 0 61 56 0 0 4
917 585
917 580
922 580
922 528
0 4 18 0 0 8320 0 0 61 130 0 4
610 558
610 695
890 695
890 649
0 3 17 0 0 8320 0 0 61 129 0 4
620 549
620 686
881 686
881 649
0 2 16 0 0 8320 0 0 61 128 0 4
629 540
629 676
872 676
872 649
1 0 15 0 0 8320 0 61 0 0 127 4
863 649
863 667
638 667
638 531
9 0 52 0 0 4096 0 61 0 0 101 2
944 649
944 799
3 5 53 0 0 4224 0 58 61 0 0 3
1023 770
899 770
899 649
3 6 54 0 0 4224 0 57 61 0 0 3
1022 737
908 737
908 649
3 7 55 0 0 4224 0 59 61 0 0 3
1023 701
917 701
917 649
3 8 56 0 0 4224 0 60 61 0 0 3
1022 668
926 668
926 649
2 0 14 0 0 4224 0 60 0 0 110 3
1071 659
1188 659
1188 557
2 0 13 0 0 8320 0 59 0 0 109 3
1072 692
1200 692
1200 548
2 0 12 0 0 8320 0 57 0 0 108 3
1071 728
1211 728
1211 539
0 2 11 0 0 4224 0 0 58 107 0 3
1220 530
1220 761
1072 761
1 0 52 0 0 0 0 58 0 0 101 2
1072 779
1102 779
1 0 52 0 0 0 0 57 0 0 101 2
1071 746
1102 746
1 0 52 0 0 0 0 59 0 0 101 2
1072 710
1102 710
1 1 52 0 0 12416 0 60 14 0 0 6
1071 677
1102 677
1102 799
290 799
290 484
144 484
1 0 37 0 0 0 0 63 0 0 116 2
1075 421
1075 369
4 0 23 0 0 8192 0 54 0 0 135 3
1320 525
1349 525
1349 283
3 0 24 0 0 8192 0 54 0 0 136 3
1320 537
1362 537
1362 277
2 0 25 0 0 8192 0 54 0 0 137 3
1320 549
1373 549
1373 271
1 0 26 0 0 8192 0 54 0 0 138 3
1320 561
1383 561
1383 265
8 15 11 0 0 0 0 54 62 0 0 4
1272 525
1253 525
1253 530
1168 530
16 7 12 0 0 0 0 62 54 0 0 4
1168 539
1271 539
1271 537
1272 537
6 17 13 0 0 0 0 54 62 0 0 4
1272 549
1271 549
1271 548
1168 548
5 18 14 0 0 0 0 54 62 0 0 4
1272 561
1253 561
1253 557
1168 557
7 0 23 0 0 8192 0 62 0 0 135 3
1104 530
1022 530
1022 283
8 0 24 0 0 8192 0 62 0 0 136 3
1104 539
1014 539
1014 277
9 0 25 0 0 0 0 62 0 0 137 3
1104 548
1005 548
1005 271
0 10 26 0 0 0 0 0 62 138 0 3
997 265
997 557
1104 557
1 0 37 0 0 0 0 64 0 0 116 2
498 431
498 369
1 0 37 0 0 12416 0 15 0 0 0 4
143 468
290 468
290 369
1478 369
8 0 23 0 0 0 0 55 0 0 135 3
742 526
772 526
772 283
7 0 24 0 0 0 0 55 0 0 136 3
742 538
785 538
785 277
6 0 25 0 0 8192 0 55 0 0 137 3
742 550
796 550
796 271
5 0 26 0 0 8192 0 55 0 0 138 3
742 562
806 562
806 265
0 1 39 0 0 4224 0 0 23 0 0 4
1480 342
254 342
254 416
146 416
0 1 27 0 0 4224 0 0 21 0 0 4
1480 330
240 330
240 382
146 382
0 1 40 0 0 4224 0 0 25 0 0 4
1481 324
232 324
232 366
146 366
0 1 41 0 0 4224 0 0 24 0 0 4
1481 318
225 318
225 349
147 349
0 1 42 0 0 4224 0 0 26 0 0 4
1481 311
218 311
218 333
146 333
0 1 43 0 0 4224 0 0 27 0 0 4
1481 305
211 305
211 315
147 315
4 15 15 0 0 0 0 55 67 0 0 4
694 526
676 526
676 531
591 531
16 3 16 0 0 0 0 67 55 0 0 3
591 540
694 540
694 538
2 17 17 0 0 0 0 55 67 0 0 3
694 550
694 549
591 549
1 18 18 0 0 0 0 55 67 0 0 4
694 562
676 562
676 558
591 558
7 0 23 0 0 8192 0 67 0 0 135 3
527 531
445 531
445 283
8 0 24 0 0 8192 0 67 0 0 136 3
527 540
437 540
437 277
9 0 25 0 0 0 0 67 0 0 137 3
527 549
428 549
428 271
0 10 26 0 0 0 0 0 67 138 0 3
420 265
420 558
527 558
8 1 23 0 0 12416 0 68 5 0 0 5
278 216
302 216
302 283
1432 283
1432 246
7 2 24 0 0 12416 0 68 5 0 0 7
278 204
308 204
308 277
1367 277
1367 278
1420 278
1420 246
6 3 25 0 0 12416 0 68 5 0 0 5
278 192
314 192
314 271
1408 271
1408 246
5 4 26 0 0 12416 0 68 5 0 0 7
278 180
319 180
319 265
1388 265
1388 266
1396 266
1396 246
19
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
1399 100 1430 129
1410 109 1418 128
1 Z
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 7
731 196 815 221
741 204 804 221
7 ALU_OUT
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
785 175 815 200
795 183 804 200
1 Z
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
784 154 814 179
794 162 803 179
1 X
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
785 130 815 155
795 138 804 155
1 B
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
784 107 814 132
794 115 803 132
1 A
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 8
7 440 100 465
17 448 89 465
8 MEMORY R
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 8
10 424 103 449
20 432 92 449
8 MEMORY W
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 4
506 144 563 169
516 152 552 169
4 DBUS
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 5
38 452 117 480
52 463 102 483
5 CLOCK
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 7
24 469 123 497
38 480 108 500
7 ADD/SUB
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
-9 405 118 430
0 411 108 428
12 DBUS=ALU_OUT
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
46 387 119 412
55 393 109 410
6 DBUS=Z
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
48 369 119 394
56 376 110 393
6 DBUS=X
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
48 353 119 378
56 359 110 376
6 DBUS=B
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 6
49 336 122 361
58 343 112 360
6 DBUS=A
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 7
42 320 122 345
50 326 113 343
7 B<-DBUS
-15 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 7
42 302 122 327
50 309 113 326
7 A<-DBUS
-27 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
47 172 77 216
54 179 69 209
1 X
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
